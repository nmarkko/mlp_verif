`include "tests/test_base.sv"
`include "tests/test_mlp_simple.sv"

