`include "sequences/axil_base_seq.sv"
`include "sequences/axis_base_seq.sv"
`include "sequences/axil_seq.sv"
`include "sequences/axis_seq.sv"
